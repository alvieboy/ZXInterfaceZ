--
--  USB Host FS controller
--
--  Copyright 2016-2020 Alvaro Lopes <alvieboy@alvie.com>
--
--  The FreeBSD license
--
--  Redistribution and use in source and binary forms, with or without
--  modification, are permitted provided that the following conditions
--  are met:
--
--  1. Redistributions of source code must retain the above copyright
--     notice, this list of conditions and the following disclaimer.
--  2. Redistributions in binary form must reproduce the above
--     copyright notice, this list of conditions and the following
--     disclaimer in the documentation and/or other materials
--     provided with the distribution.
--
--  THIS SOFTWARE IS PROVIDED BY THE AUTHOR ``AS IS'' AND ANY
--  EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
--  THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
--  PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
--  ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
--  INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
--  (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
--  OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
--  HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
--  STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
--  ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
--  ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--
--


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;
library work;
use work.usbpkg.all;
use work.ahbpkg.all;
-- synopsys translate_off
use work.txt_util.all;
-- synopsys translate_on

ENTITY usbhostctrl IS
  PORT (
    usbclk_i    : in std_logic;
    ausbrst_i   : in std_logic;

    -- Comms to external world
    ahb_m2s_i   : in AHB_M2S;
    ahb_s2m_o   : out AHB_S2M;


    clk_i       : in std_logic;
    arst_i      : in std_logic;
    int_o       : out std_logic; -- sync to clk_i
    int_async_o : out std_logic; -- sync to usb clock
    -- Interface to transceiver
    softcon_o   : out std_logic;
    noe_o       : out std_logic;
    speed_o     : out std_logic;
    vpo_o       : out std_logic;
    vmo_o       : out std_logic;
    mode_o      : out std_logic;
    suspend_o   : out std_logic;

    rcv_i       : in std_logic;
    vp_i        : in  std_logic;
    vm_i        : in  std_logic;
    pwren_o     : out std_logic;
    pwrflt_i    : in std_logic;
    dbg_o       : out std_logic_vector(7 downto 0)
  );
END entity usbhostctrl;

ARCHITECTURE rtl OF usbhostctrl is

  SIGNAL  Phy_DataIn     : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL  Phy_DataOut    : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL  Phy_Linestate  : STD_LOGIC_VECTOR(1 DOWNTO 0);
  SIGNAL  Phy_Opmode     : STD_LOGIC_VECTOR(1 DOWNTO 0);
  SIGNAL  Phy_RxActive   : STD_LOGIC;
  SIGNAL  Phy_RxError    : STD_LOGIC;
  SIGNAL  Phy_RxValid    : STD_LOGIC;
  SIGNAL  Phy_Termselect : STD_LOGIC := 'L';
  SIGNAL  Phy_TxReady    : STD_LOGIC;
  SIGNAL  Phy_TxValid    : STD_LOGIC;
  SIGNAL  Phy_XcvrSelect : STD_LOGIC := 'L';
  SIGNAL  usb_rst_phy    : STD_LOGIC;
  SIGNAL  usb_rst_slv    : STD_LOGIC;

  signal rstinv         : std_logic;
  signal tx_mode_s      : std_logic := '1';
  signal rst_event_q    : std_logic;
  signal rst_event      : std_logic;
  signal noe_s          : std_logic;

  signal rd_s           : std_logic;
  signal wr_s           : std_logic;
  signal addr_s         : std_logic_vector(11 downto 0);
  signal dat_in_s       : std_logic_vector(7 downto 0);
  signal dat_out_s      : std_logic_vector(7 downto 0);




  signal dbg_rx_data_done_s : std_logic;
  signal dbg_trans_state_s  : std_logic_vector(4 downto 0);
  signal cnt_ack_s       : std_logic_vector(7 downto 0);
  signal cnt_nack_s      : std_logic_vector(7 downto 0);
  signal cnt_babble_s    : std_logic_vector(7 downto 0);
  signal cnt_stall_s     : std_logic_vector(7 downto 0);
  signal cnt_crcerror_s  : std_logic_vector(7 downto 0);
  signal cnt_timeout_s   : std_logic_vector(7 downto 0);
  signal cnt_errorpid_s  : std_logic_vector(7 downto 0);
  signal cnt_cplt_s      : std_logic_vector(7 downto 0);

  constant C_SOF_TIMEOUT: natural   := altsim(48000, 4800*2); -- 1ms, 100us
  constant C_ATTACH_DELAY: natural  := altsim(480000, 4);-- 48000; -- 10 ms
  constant C_NUM_CHANNELS: natural  := 8;
  constant C_RESET_DELAY: natural   := altsim(48000*50,500); -- 50 ms
  constant C_RESET_DELAY_AFTER: natural   := altsim(480, 48); -- 10 us
  constant C_INTERRUPT_HOLDOFF : natural := altsim(4800*5, 480); -- 500us / 10us

  signal dbg_chan_interrupt_s : std_logic_vector(C_NUM_CHANNELS-1 downto 0);

  type host_state_type is (
    DETACHED,
    ATTACHED,
    IDLE,
    RESET1,
    RESET2,
    --SUSPEND,
    --RESUME,
    WAIT_SOF,
    IN1,
    OUT1,
    SOF1,
    SETUP1
  );

  type status_reg_type is record
    fulllowspeed    : std_logic; -- '1': FS, '0': LS
    poweron         : std_logic;
    reset           : std_logic;
    suspend         : std_logic;
    overcurrent     : std_logic;
    --connectdetect   : std_logic;
    connected       : std_logic;
  end record;

  type interrupt_reg_type is record
    overcurrent     : std_logic; -- Interrupt on overcurrent
    connectdetect   : std_logic; -- Interrupt on connect event
    disconnectdetect: std_logic; -- Interrupt on disconnect event
    ginten          : std_logic; -- Global USB interrupt enable
  end record;

  constant C_EP_TYPE_INTERRUPT: std_logic_vector(1 downto 0) := "11";

  type channel_conf_reg_type is record
    enabled         : std_logic;
    oddframe        : std_logic;
    lowspeed        : std_logic;
    direction       : std_logic;
    epnum           : std_logic_vector(3 downto 0);
    address         : std_logic_vector(6 downto 0);
    eptype          : std_logic_vector(1 downto 0); -- 00: Control
                                                    -- 01: Isochronous
                                                    -- 10: Bulk
                                                    -- 11: Interrupt

    maxsize         : std_logic_vector(5 downto 0); -- Max 64 bytes.
    interval        : std_logic_vector(7 downto 0); -- for interrupt endpoints
  end record;

  constant C_RESET_CHANNEL_CONF: channel_conf_reg_type := (
    '0',
    'X',
    'X',
    'X',
    (others => 'X'),
    (others => 'X'),
    (others => 'X'),
    (others => 'X'),
    (others => '0')
  );

  type channel_trans_reg_type is record
    dpid            : std_logic_vector(1 downto 0);  -- Data PID.;
                                                     -- 11: setup
                                                     -- 00: IN
                                                     -- 01: OUT
    cnt             : std_logic; -- Limited to 1 packet.
    seq             : std_logic;
    size            : unsigned(6 downto 0);
    epaddr          : unsigned(9 downto 0);
    retries         : unsigned(1 downto 0);
    intervalcnt     : unsigned(7 downto 0); -- for interrupt endpoints
    issued          : std_logic;
  end record;

  constant C_RESET_TRANS: channel_trans_reg_type := (
    (others => 'X'),
    'X',
    'X',
    (others => 'X'),
    (others => 'X'),
    (others => 'X'),
    (others => 'X'),
    'X'
  );

  type channel_interrupt_conf_reg_type is record
    datatogglerror  : std_logic;
    crcerror        : std_logic;
    babble          : std_logic;
    transerror      : std_logic; -- Timeout
                                 -- Bit stuff error
                                 -- False EOP
    ack             : std_logic;
    nack            : std_logic;
    stall           : std_logic;
    cplt            : std_logic; -- Completed
  end record;

  constant C_RESET_INTERRUPT_CONF: channel_interrupt_conf_reg_type := ( others => 'X' );
  constant C_RESET_INTERRUPT_PEND: channel_interrupt_conf_reg_type := ( others => '0' );


  type channel_type is record
    conf      : channel_conf_reg_type;
    trans     : channel_trans_reg_type;
    intconf   : channel_interrupt_conf_reg_type;
    intpend   : channel_interrupt_conf_reg_type;
  end record;

  type channels_type is array (0 to C_NUM_CHANNELS-1) of channel_type;

  type regs_type is record
    host_state      : host_state_type;
    sr              : status_reg_type;
    intconfr        : interrupt_reg_type;
    intpendr        : interrupt_reg_type;
    speed           : std_logic;
    attach_count    : natural range 0 to C_ATTACH_DELAY - 1;
    sof_count       : natural range 0 to C_SOF_TIMEOUT - 1;
    frame           : unsigned(10 downto 0);
    channel         : natural range 0 to C_NUM_CHANNELS -1;
    reset_delay     : natural range 0 to C_RESET_DELAY-1;
    ch              : channels_type;
    int_holdoff     : natural range 0 to C_INTERRUPT_HOLDOFF-1;
  end record;

  signal r                    : regs_type := (
    DETACHED,
    ( others => 'X'),
    ( others => 'X'),
    ( others => 'X'),
    'X',
    C_ATTACH_DELAY-1,
    C_SOF_TIMEOUT-1,
    ( others => 'X'),
    0,
    C_RESET_DELAY-1,
    ( others => ( C_RESET_CHANNEL_CONF,
      C_RESET_TRANS,
      C_RESET_INTERRUPT_CONF,
      C_RESET_INTERRUPT_PEND
      )
    ),
    C_INTERRUPT_HOLDOFF-1
  );
  --signal frame_crc5_s         : std_logic_vector(4 downto 0);

  signal statusreg_s          : std_logic_vector(7 downto 0);
  --signal intconfreg_s         : std_logic_vector(7 downto 0);
  signal intpendreg_s         : std_logic_vector(7 downto 0);

  --signal write_data_s         : std_logic_vector(7 downto 0);
  --signal write_address_s      : std_logic_vector(10 downto 0);


  signal vpo_s, vmo_s: std_logic;



  signal address_ep_crc_in_s: std_logic_vector(10 downto 0);
  signal address_ep_crc_out_s: std_logic_vector(4 downto 0);

  signal debug_ch:  channel_type;

  -- Epmem
  signal epmem_read_en_s    : std_logic;
  signal epmem_write_en_s   : std_logic;
  signal epmem_addr_s       : std_logic_vector(9 downto 0);
  signal epmem_data_in_s    : std_logic_vector(7 downto 0);
  signal epmem_data_out_s   : std_logic_vector(7 downto 0);
  signal hep_dat_s          : std_logic_vector(7 downto 0);
  signal hep_rd_s   : std_logic;
  signal hep_wr_s   : std_logic;



  signal int_s                : std_logic;
  signal int_sync_s           : std_logic;
  signal read_data_s          : std_logic_vector(7 downto 0);

  signal trans_addr_s       : std_logic_vector(6 downto 0);
  signal trans_dsize_s      : std_logic_vector(6 downto 0);
  signal trans_dsize_read_s : std_logic_vector(6 downto 0);
  signal trans_daddr_s      : std_logic_vector(9 downto 0);
  signal trans_ep_s         : std_logic_vector(3 downto 0);
  signal trans_status_s     : usb_transaction_status_type;
  signal trans_pid_s        : std_logic_vector(3 downto 0);
  signal trans_strobe_s     : std_logic;
  signal trans_data_seq_s   : std_logic;
  signal trans_seq_valid_s  : std_logic;
  signal trans_speed_s      : std_logic;
  signal phy_txactive_s     : std_logic;
  signal fs_ce_s            : std_logic;
	signal dbg_fs_ce_r		: std_logic;
  signal read_data_r        : std_logic_vector(7 downto 0);
BEGIN

  rstinv      <= not ausbrst_i;
  suspend_o   <= '0';

  statusreg_s <= '0' &
    r.sr.fulllowspeed & 
    r.sr.poweron      & 
    r.sr.reset        &
    '0' & --r.sr.suspend       &
    r.sr.overcurrent   &
    '0' &
    r.sr.connected;

  --intconfreg_s <= r.intconfr.ginten & "0000" & r.intconfr.overcurrent & r.intconfr.connectdetect & r.intconfr.disconnectdetect;
  intpendreg_s <= "00000" & r.intpendr.overcurrent & r.intpendr.connectdetect & r.intpendr.disconnectdetect;


  
  usb_phy_inst : ENTITY work.usb_phy       --Open Cores USB Phy, designed by Rudolf Usselmanns
  GENERIC MAP (
    usb_rst_det      => TRUE,
    CLOCK            => "48"
  )
  PORT MAP (
    clk              => usbclk_i,       -- i
    rst              => rstinv,         -- i
    phy_tx_mode      => tx_mode_s,      -- i
    usb_rst          => usb_rst_phy,    -- o
    XcvrSelect_i     => Phy_XcvrSelect,--r.speed,        -- i
    HostXcvrSelect_i => r.speed,
    fs_ce_o          => fs_ce_s,
    txdp             => vpo_s,          -- o
    txdn             => vmo_s,          -- o
    txoe             => noe_s,          -- o
    rxd              => rcv_i,          -- i
    rxdp             => vp_i,           -- i
    rxdn             => vm_i,           -- i
    DataOut_i        => Phy_DataOut,    -- i (7 downto 0);
    TxValid_i        => Phy_TxValid,    -- i
    TxReady_o        => Phy_TxReady,    -- o
    DataIn_o         => Phy_DataIn,     -- o (7 downto 0);
    RxValid_o        => Phy_RxValid,    -- o
    RxActive_o       => Phy_RxActive,   -- o
    RxError_o        => Phy_RxError,    -- o
    LineState_o      => Phy_LineState   -- o (1 downto 0). (0) is P, (1) is N
  );

  phy_txactive_s <= not noe_s;

  mainp: process(usbclk_i, ausbrst_i, r, Phy_Linestate, dat_in_s, addr_s, rd_s, wr_s, statusreg_s, intpendreg_s,
    usb_rst_phy, trans_status_s, trans_dsize_read_s, pwrflt_i)
    variable w  : regs_type;
    variable ch : channel_type;
    variable wch_u : unsigned(2 downto 0);
    variable wch : natural;
    variable channel_handled: boolean;
    variable can_issue_request: boolean;
    variable interrupt_v: std_logic_vector(C_NUM_CHANNELS-1 downto 0);
  begin
    w := r;
    tx_mode_s       <= '1';
    -- Optimizations
    trans_pid_s     <= (others => 'X');
    trans_strobe_s  <= '0';
    trans_addr_s    <= (others => 'X');
    trans_dsize_s   <= (others => 'X');
    trans_daddr_s   <= (others => 'X');
    trans_ep_s      <= (others => 'X');
    trans_data_seq_s<='X';
    trans_speed_s   <= 'X';--not r.ch(r.channel).trans.lowspeed;
    --trans_addr_s    <= (others => 'X');
    read_data_s     <= (others => '0');

    -- End optimizations
    if r.sof_count=0 then
      w.sof_count         := C_SOF_TIMEOUT - 1;
      w.frame             := r.frame + 1;
    else
      w.sof_count         := r.sof_count - 1;
    end if;

    chint: for i in 0 to C_NUM_CHANNELS-1 loop
      interrupt_v(i) := '0';
      if  r.ch(i).intpend.datatogglerror = '1' or
          r.ch(i).intpend.crcerror       = '1' or
          r.ch(i).intpend.babble         = '1' or
          r.ch(i).intpend.transerror     = '1' or
          r.ch(i).intpend.ack            = '1' or
          r.ch(i).intpend.nack           = '1' or
          r.ch(i).intpend.stall          = '1' or
          r.ch(i).intpend.cplt           = '1'
         then
        interrupt_v(i) := '1';
      end if;
    end loop;

    --if r.int_holdoff=0 then
      int_s <= (or_reduce(interrupt_v) or r.intpendr.connectdetect or r.intpendr.overcurrent
        or r.intpendr.disconnectdetect ) and r.intconfr.ginten;
    dbg_chan_interrupt_s <= interrupt_v;
    --else
    --  int_s <= '0';
    --  w.int_holdoff := r.int_holdoff - 1;
    --end if;

    -- Process writes coming from SPI
    if wr_s='1' then
      if addr_s(10 downto 7) = "0000" then
        case addr_s(6 downto 0) is
          when "0000000" =>
            w.sr.poweron               := dat_in_s(5);
            if dat_in_s(4)='1' then w.sr.reset := '1'; end if;

          when "0000010" =>  -- Interrupt conf reg
            w.intconfr.ginten         := dat_in_s(7);
            w.intconfr.disconnectdetect  := dat_in_s(0);
            w.intconfr.connectdetect  := dat_in_s(1);
            w.intconfr.overcurrent    := dat_in_s(2);
          when "0000011" =>
            -- Interrupt clear/ack
            if dat_in_s(0)='1' then w.intpendr.disconnectdetect := '0'; end if;
            if dat_in_s(1)='1' then w.intpendr.connectdetect := '0'; end if;
            if dat_in_s(2)='1' then w.intpendr.overcurrent   := '0'; end if;
            if dat_in_s(7)='1' then w.int_holdoff:=C_INTERRUPT_HOLDOFF-1; end if;
    
          when others =>
        end case;
      elsif addr_s(10 downto 7) = "0001" then
          wch_u := unsigned(addr_s(6 downto 4));
          wch := to_integer(wch_u);
          case addr_s(3 downto 0) is
            when "0000" =>
              w.ch(wch).conf.eptype    := dat_in_s(7 downto 6);
              w.ch(wch).conf.maxsize   := dat_in_s(5 downto 0);
            when "0001" =>
              --w.ch(wch).conf.oddframe  := dat_in_s(7);
              w.ch(wch).conf.direction := dat_in_s(7);
              w.ch(wch).conf.lowspeed  := dat_in_s(6);
              w.ch(wch).conf.epnum     := dat_in_s(3 downto 0);

            when "0010" =>
              w.ch(wch).conf.enabled   := dat_in_s(7);
              w.ch(wch).conf.address   := dat_in_s(6 downto 0);
            when "0011" => -- Interrupt configuration
              w.ch(wch).intconf.datatogglerror  := dat_in_s(7);
              w.ch(wch).intconf.crcerror    := dat_in_s(6);
              w.ch(wch).intconf.babble          := dat_in_s(5);
              w.ch(wch).intconf.transerror      := dat_in_s(4);
              w.ch(wch).intconf.ack             := dat_in_s(3);
              w.ch(wch).intconf.nack            := dat_in_s(2);
              w.ch(wch).intconf.stall           := dat_in_s(1);
              w.ch(wch).intconf.cplt            := dat_in_s(0);
            when "0100" => -- Interrupt clear
              if dat_in_s(7)='1' then w.ch(wch).intpend.datatogglerror  := '0'; end if;
              if dat_in_s(6)='1' then w.ch(wch).intpend.crcerror        := '0'; end if;
              if dat_in_s(5)='1' then w.ch(wch).intpend.babble          := '0'; end if;
              if dat_in_s(4)='1' then w.ch(wch).intpend.transerror      := '0'; end if;
              if dat_in_s(3)='1' then w.ch(wch).intpend.ack             := '0'; end if;
              if dat_in_s(2)='1' then w.ch(wch).intpend.nack            := '0'; end if;
              if dat_in_s(1)='1' then w.ch(wch).intpend.stall           := '0'; end if;
              if dat_in_s(0)='1' then w.ch(wch).intpend.cplt            := '0'; end if;

            when "0101" =>
              w.ch(wch).conf.interval       := dat_in_s;
              w.ch(wch).trans.intervalcnt   := unsigned(dat_in_s); -- restart counter.
            when "1000" =>
              w.ch(wch).trans.dpid    := dat_in_s(1 downto 0);
              w.ch(wch).trans.seq     := dat_in_s(2);
              w.ch(wch).trans.epaddr(9 downto 8)  := unsigned(dat_in_s(4 downto 3));
              w.ch(wch).trans.retries := unsigned(dat_in_s(6 downto 5));

            when "1001" => -- Transaction
              w.ch(wch).trans.epaddr(7 downto 0)   := unsigned(dat_in_s);

            when "1010" => -- Transaction
              w.ch(wch).trans.size := unsigned(dat_in_s(6 downto 0));
              w.ch(wch).trans.cnt  := dat_in_s(7);
            when others =>
          end case;
      end if;
    end if;

    -- read data
    if not is_x(addr_s) and rd_s='1' then

      if addr_s(10 downto 7) = "0000" then
        case addr_s(6 downto 0) is
          when "0000000" =>
            read_data_s <= statusreg_s;
          when "0000001" =>
            -- channel interrupt pending reg
            read_data_s <= intpendreg_s;
          when "0000010" =>
            --  interrupt status reg
            read_data_s <= interrupt_v;

          when "0000011" =>

            case trans_status_s is
              when IDLE       =>  read_data_s <= x"00";
              when BUSY       =>  read_data_s <= x"01";
              when TIMEOUT    =>  read_data_s <= x"02";
              when BABBLE     =>  read_data_s <= x"03";
              when ACK        =>  read_data_s <= x"04";
              when NACK       =>  read_data_s <= x"05";
              when STALL      =>  read_data_s <= x"06";
              when CRCERROR   =>  read_data_s <= x"07";
              when COMPLETED  =>  read_data_s <= x"08";
              when others     =>  read_data_s <= x"0F";
            end case;

          when "0000100" =>
            case r.host_state is
              when DETACHED   =>  read_data_s <= x"00";
              when ATTACHED   =>  read_data_s <= x"01";
              when IDLE       =>  read_data_s <= x"02";
              when RESET1     =>  read_data_s <= x"03";
              when RESET2     =>  read_data_s <= x"04";
              when WAIT_SOF   =>  read_data_s <= x"05";
              when IN1        =>  read_data_s <= x"06";
              when OUT1       =>  read_data_s <= x"07";
              when SETUP1     =>  read_data_s <= x"08";
              when SOF1       =>  read_data_s <= x"09";
              when others     =>  read_data_s <= x"0F";
            end case;
          when "0000101" =>

            read_data_s <= "000" & dbg_trans_state_s ;

          when "0000110" =>
              read_data_s <= cnt_ack_s;
          when "0000111" =>
              read_data_s <= cnt_nack_s;
          when "0001000" =>
              read_data_s <= cnt_babble_s;
          when "0001001" =>
              read_data_s <= cnt_stall_s;
          when "0001010" =>
              read_data_s <= cnt_crcerror_s;
          when "0001011" =>
              read_data_s <= cnt_timeout_s;
          when "0001100" =>
              read_data_s <= cnt_errorpid_s;
          when "0001101" =>
              read_data_s <= cnt_cplt_s;
          when others =>
            read_data_s <= (others =>'X');
        end case;

      elsif addr_s(10 downto 7) = "0001" then
        wch_u := unsigned(addr_s(6 downto 4));
        wch := to_integer(wch_u);
        case addr_s(3 downto 0) is
          when "0000" =>
            read_data_s(7 downto 6) <= r.ch(wch).conf.eptype;
            read_data_s(5 downto 0) <= r.ch(wch).conf.maxsize;
          when "0001" =>
            --read_data_s(7)          <= r.ch(wch).conf.oddframe;
            read_data_s(6)          <= r.ch(wch).conf.lowspeed;
            read_data_s(7)          <= r.ch(wch).conf.direction;
            read_data_s(3 downto 0) <= r.ch(wch).conf.epnum;
          --
          when "0010" =>
            read_data_s(7)          <= r.ch(wch).conf.enabled;
            read_data_s(6 downto 0) <= r.ch(wch).conf.address;
          when "0011" => -- Interrupt configuration
            read_data_s(7)          <= r.ch(wch).intconf.datatogglerror;
            read_data_s(6)          <= r.ch(wch).intconf.crcerror;
            read_data_s(5)          <= r.ch(wch).intconf.babble;
            read_data_s(4)          <= r.ch(wch).intconf.transerror;
            read_data_s(3)          <= r.ch(wch).intconf.ack;
            read_data_s(2)          <= r.ch(wch).intconf.nack;
            read_data_s(1)          <= r.ch(wch).intconf.stall;
            read_data_s(0)          <= r.ch(wch).intconf.cplt;
          when "0100" => -- Interrupt read
            read_data_s(7)          <= r.ch(wch).intpend.datatogglerror;
            read_data_s(6)          <= r.ch(wch).intpend.crcerror;
            read_data_s(5)          <= r.ch(wch).intpend.babble;
            read_data_s(4)          <= r.ch(wch).intpend.transerror;
            read_data_s(3)          <= r.ch(wch).intpend.ack;
            read_data_s(2)          <= r.ch(wch).intpend.nack;
            read_data_s(1)          <= r.ch(wch).intpend.stall;
            read_data_s(0)          <= r.ch(wch).intpend.cplt;
          when "0101" =>
            read_data_s             <= r.ch(wch).conf.interval;
          when "1000" =>
            read_data_s(1 downto 0) <= r.ch(wch).trans.dpid;
            read_data_s(2)          <= r.ch(wch).trans.seq;
            read_data_s(4 downto 3) <= std_logic_vector(r.ch(wch).trans.epaddr(9 downto 8));
            read_data_s(6 downto 5) <= std_logic_vector(r.ch(wch).trans.retries);
          when "1001" => -- Transaction
            read_data_s             <= std_logic_vector(r.ch(wch).trans.epaddr(7 downto 0));
          when "1010" => -- Transaction
            read_data_s(6 downto 0) <= std_logic_vector(r.ch(wch).trans.size);
            read_data_s(7)          <= r.ch(wch).trans.cnt;
          when others =>
            read_data_s <= (others => 'X');
          end case;
      else
        read_data_s <= (others => 'X');
      end if;
    else
      read_data_s <= (others => 'X');
    end if;

    ch := r.ch( r.channel );
    debug_ch <= ch;

    case r.host_state is
      when DETACHED =>
        if not is_x(Phy_Linestate) and ( Phy_Linestate="01" or Phy_Linestate="10" ) then
          if r.sr.poweron='1' then
          if r.attach_count=0 then
            w.sr.fulllowspeed   := Phy_Linestate(0); -- Set speed according to USB+ pullup
            w.speed := Phy_Linestate(0); -- Set speed according to USB+ pullup
            w.host_state        := ATTACHED;
            --w.sr.connectdetect  :='1';
            -- synthesis translate_off
            report "DEVICE ATTACHED";-- severity failure;
            -- synthesis translate_on
            w.sr.connected      :='1';
            if r.intconfr.connectdetect='1' then
              w.intpendr.connectdetect:='1';
            end if;
            w.sof_count         := C_SOF_TIMEOUT - 1;
          else
            w.attach_count      := r.attach_count - 1;
          end if;
          end if;
        else
          w.attach_count        := C_ATTACH_DELAY - 1;
          --w.sr.connectdetect    :='0';
          w.sr.connected        :='0';
        end if;

      when ATTACHED | IDLE =>

        channel_handled   := false;
        can_issue_request := false;
        --
        -- sync   pid  +packet  crc
        --
        -- 8    + 8    512[s]  + 16    528 bits, 105 blocks of 5 bits. 3 extra bits. 633 bits MAX. 649 bits incl. sync+pid
        -- 8    + 8    64[s]   + 16    80 bits, 96 bits MAX. 112 bits incl. sync+pid     4600.

        --34 bits time for ack/nack . 38 bits for token.

        -- Counter starts at 4799

        if ch.conf.lowspeed='0' then -- High speed (64 bytes)
          if r.sof_count > ((649+34+38)*4) then
            can_issue_request := true;
          end if;
        else                      -- Low speed (8 bytes)
          if r.sof_count > ((112+34+38)*4*8) then -- TBD: this is wrong!
            can_issue_request := true;
          end if;
        end if;
        -- synthesis translate_off
        --  if r.sof_count > 100 then
        --    can_issue_request := true;
        --  end if;
        -- synthesis translate_on

        if ch.conf.enabled='1' then
          -- synopsys translate_off
          if rising_edge(usbclk_i) then
            --report "Channel "&str(r.channel)&" enabled";
          end if;
          -- synopsys translate_on

          if ch.conf.eptype = C_EP_TYPE_INTERRUPT and (ch.trans.intervalcnt/=0 or ch.trans.issued='1')then
            can_issue_request := false;
          end if;

          if ch.trans.cnt/='0' and can_issue_request then
            if ch.trans.dpid="11" then
              report "Got setup request";
              w.host_state := SETUP1;
              channel_handled := true;
            elsif ch.trans.dpid="00" and ch.trans.issued='0' then    -- Do not retry IN ad infinitum
              w.host_state := IN1;
              channel_handled := true;
            elsif ch.trans.dpid="01" then
              w.host_state := OUT1;
              channel_handled := true;
            end if;
          end if;
        end if;

        if r.sr.reset='1' then
          w.host_state := RESET1;
          w.reset_delay := C_RESET_DELAY -1;
        end if;

        if not channel_handled then
          if r.channel /= C_NUM_CHANNELS-1 then
            w.channel := r.channel + 1;
          else
            w.channel := 0;
            if not can_issue_request then
              w.host_state := WAIT_SOF;
            end if;
          end if;
        end if;

        if r.sr.poweron='0' then
          w.host_state := DETACHED;
        end if;

      when WAIT_SOF =>
        if r.sof_count=0 then
          w.host_state := SOF1;
        end if;
        if r.sr.reset='1' then
          w.host_state := RESET1;
          w.reset_delay := C_RESET_DELAY -1;
        end if;

        if r.sr.poweron='0' then
          w.host_state := DETACHED;
        end if;
          if usb_rst_phy='1' then
          -- Disconnected???
            if r.intconfr.disconnectdetect='1' then
              w.intpendr.disconnectdetect := '1';
            end if;
            w.sr.connected := '0';
            w.host_state := DETACHED;
          end if;


      when SOF1 =>
        trans_pid_s     <= USBF_T_PID_SOF;
        trans_strobe_s  <= '1';
        trans_speed_s   <= r.sr.fulllowspeed;

        if trans_status_s=COMPLETED then
          -- For all interrupt EPs, decrease counters
          ie: for i in 0 to C_NUM_CHANNELS-1 loop
            w.ch(i).trans.issued := '0';

            --if r.ch(i).conf.eptype = C_EP_TYPE_INTERRUPT then
              if r.ch(i).trans.intervalcnt=0 then
                w.ch(i).trans.intervalcnt := unsigned(r.ch(i).conf.interval);
              else
                w.ch(i).trans.intervalcnt := r.ch(i).trans.intervalcnt - 1;
              end if;
            --end if;
          end loop;

          w.host_state := IDLE;
        end if;

      when SETUP1 =>
        trans_pid_s       <= USBF_T_PID_SETUP;
        trans_strobe_s    <= '1';

        trans_daddr_s     <= std_logic_vector(r.ch(r.channel).trans.epaddr);
        trans_dsize_s     <= std_logic_vector(r.ch(r.channel).trans.size);
        trans_ep_s        <= r.ch(r.channel).conf.epnum;
        trans_addr_s      <= r.ch(r.channel).conf.address;
        trans_data_seq_s  <= r.ch(r.channel).trans.seq;
        trans_speed_s     <= not r.ch(r.channel).conf.lowspeed;

        case trans_status_s is
          when ACK =>
            -- synthesis translate_off
            if rising_edge(usbclk_i) then report "Got ACK for SETUP"; end if;
            -- synthesis translate_on

            w.ch(r.channel).trans.cnt   := '0';
            w.ch(r.channel).intpend.ack := '1';
            w.ch(r.channel).intpend.cplt:= '1';
            w.host_state := IDLE;
          when NACK =>
            -- Keep trying...
            w.host_state := IDLE;

          when STALL =>
            w.ch(r.channel).intpend.stall := '1';
            w.ch(r.channel).trans.cnt   := '0';
            w.host_state := IDLE;

          when IDLE | BUSY =>
            -- Stay here.
          when others =>
            w.ch(r.channel).trans.cnt   := '0';
            w.ch(r.channel).intpend.transerror := '1';
            w.host_state := IDLE;
        end case;


      when IN1 =>
        trans_pid_s     <= USBF_T_PID_IN;
        trans_strobe_s  <= '1';

        trans_daddr_s   <= std_logic_vector(r.ch(r.channel).trans.epaddr);
        trans_dsize_s   <= std_logic_vector(r.ch(r.channel).trans.size);
        trans_ep_s      <= r.ch(r.channel).conf.epnum;
        trans_addr_s    <= r.ch(r.channel).conf.address;
        trans_data_seq_s  <= r.ch(r.channel).trans.seq;
        trans_speed_s     <= not r.ch(r.channel).conf.lowspeed;
        case trans_status_s is
          when COMPLETED =>
            w.ch(r.channel).trans.cnt    := '0';
            w.ch(r.channel).intpend.cplt := '1';
            if trans_seq_valid_s='0' then
              w.ch(r.channel).intpend.datatogglerror := '1';
            end if;
            --w.ch(r.channel).intpend.ack  := '1';

            -- TODO: check data sequence!!!

            -- synthesis translate_off
            if rising_edge(usbclk_i) then report "IN completed, len " & hstr(trans_dsize_read_s); end if;
            -- synthesis translate_on
            w.host_state := IDLE;
            w.ch(r.channel).trans.size := unsigned(trans_dsize_read_s);
          when NACK =>
            -- Keep trying...
            w.ch(r.channel).trans.issued := '1';
            -- synthesis translate_off
            if rising_edge(usbclk_i) then report "IN NAK" & hstr(trans_dsize_read_s); end if;
            -- synthesis translate_on
            w.host_state := IDLE;

          when IDLE | BUSY =>

          when TIMEOUT | CRCERROR =>
            -- Retry
            if r.ch(r.channel).trans.retries="00" then
              if trans_status_s=TIMEOUT then
                w.ch(r.channel).intpend.transerror  := '1';
              else
                w.ch(r.channel).intpend.crcerror    := '1';
              end if;
              w.ch(r.channel).trans.cnt   := '0';
            else
              w.ch(r.channel).trans.retries := r.ch(r.channel).trans.retries - 1;
            end if;
            w.host_state := IDLE;

          when BABBLE =>
            w.ch(r.channel).intpend.stall := '1';
            w.ch(r.channel).trans.cnt   := '0';
            w.host_state := IDLE;

          when STALL =>
            w.ch(r.channel).intpend.stall := '1';
            w.ch(r.channel).trans.cnt   := '0';
            w.host_state := IDLE;

          when others =>
            -- synthesis translate_off
            if rising_edge(usbclk_i) then report "Unknown state " & hstr(trans_dsize_read_s); end if;
            -- synthesis translate_on

            w.ch(r.channel).intpend.transerror := '1';
            w.ch(r.channel).trans.cnt   := '0';
            w.host_state := IDLE;
        end case;

      when OUT1 =>
        trans_pid_s     <= USBF_T_PID_OUT;
        trans_strobe_s  <= '1';

        trans_daddr_s     <= std_logic_vector(r.ch(r.channel).trans.epaddr);
        trans_dsize_s     <= std_logic_vector(r.ch(r.channel).trans.size);
        trans_ep_s        <= r.ch(r.channel).conf.epnum;
        trans_addr_s      <= r.ch(r.channel).conf.address;
        trans_data_seq_s  <= r.ch(r.channel).trans.seq;
        trans_speed_s     <= not r.ch(r.channel).conf.lowspeed;

        case trans_status_s is
          when COMPLETED  | ACK=>
            w.ch(r.channel).trans.cnt    := '0';
            w.ch(r.channel).intpend.cplt := '1';
            w.ch(r.channel).intpend.ack  := '1';

            w.ch(r.channel).trans.seq    := not r.ch(r.channel).trans.seq;
            -- synthesis translate_off
            if rising_edge(usbclk_i) then report "OUT completed, len " & hstr(trans_dsize_read_s); end if;
            -- synthesis translate_on
            w.host_state := IDLE;
            w.ch(r.channel).trans.size := unsigned(trans_dsize_read_s);
          when NACK =>
            -- Keep trying...
            -- synthesis translate_off
            if rising_edge(usbclk_i) then report "OUT NAK" & hstr(trans_dsize_read_s); end if;
            -- synthesis translate_on
            w.host_state := IDLE;

          when STALL =>
            w.ch(r.channel).intpend.stall := '1';
            w.ch(r.channel).trans.cnt   := '0';
            w.host_state := IDLE;
          when IDLE | BUSY =>

          when TIMEOUT =>
            w.ch(r.channel).trans.cnt   := '0';
            w.ch(r.channel).intpend.transerror := '1';
            w.host_state := IDLE;

          when CRCERROR =>
            w.ch(r.channel).trans.cnt   := '0';
            w.ch(r.channel).intpend.crcerror := '1';
            w.host_state := IDLE;

          when others =>
                      -- synthesis translate_off
            if rising_edge(usbclk_i) then report "Unknown state " & hstr(trans_dsize_read_s); end if;
            -- synthesis translate_on

            w.ch(r.channel).trans.cnt   := '0';
            w.ch(r.channel).intpend.transerror := '1';
            w.host_state := IDLE;
        end case;


      when RESET1 =>
        tx_mode_s <= '0'; -- Single-ended
        --Phy_DataOut <= "10101010";
        --Phy_TxValid <= '1';
        if r.reset_delay = 0 then
          w.reset_delay := C_RESET_DELAY_AFTER;
          w.host_state := RESET2;
        else
          w.reset_delay := r.reset_delay-1;
        end if;

      when RESET2 =>
        if r.reset_delay = 0 then
          w.sr.reset := '0';
          w.host_state := IDLE;
        else
          w.reset_delay := r.reset_delay-1;
        end if;

      when others =>
        report "INVALID STATE";

    end case;


    if usb_rst_phy='1' and tx_mode_s='1' then
      -- Disconnected???
      --w.sr.connectdetect := '1';
      --if r.intconfr.disconnectdetect='1' then
      --  w.intpendr.disconnectdetect := '1';
      --end if;

      --w.sr.connected := '0';
      --w.host_state := DETACHED;
    end if;


    w.sr.overcurrent := not pwrflt_i;

    if pwrflt_i='0' and r.intconfr.overcurrent='1' then
      w.intpendr.overcurrent:='1';
    end if;

                             
    if ausbrst_i='1' then
      r.host_state        <= DETACHED;
      r.frame             <= (others => '0');--"10100010101";
      r.sof_count         <= C_SOF_TIMEOUT - 1;
      r.attach_count      <= C_ATTACH_DELAY - 1;
      r.channel           <= 0;
      r.sr.poweron        <= '0';
      r.sr.overcurrent    <= '0';
      r.sr.fulllowspeed   <= '0';
      r.sr.connected      <= '0';
      r.sr.reset          <= '0';
      r.sr.suspend        <= '0';
      r.speed             <= 'X';
      r.intpendr.connectdetect <= '0';
      r.intpendr.disconnectdetect <= '0';
      r.intpendr.overcurrent   <= '0';
      r.intconfr.ginten        <= '0';
      r.intconfr.connectdetect <= '0';
      r.intconfr.disconnectdetect <= '0';
      r.intconfr.overcurrent   <= '0';
      r.int_holdoff            <= C_INTERRUPT_HOLDOFF-1;
      r.reset_delay       <= C_RESET_DELAY-1;

      chc: for i in 0 to C_NUM_CHANNELS-1 loop
        r.ch(i).conf.enabled      <= '0';
        r.ch(i).conf.direction    <= 'X';
        r.ch(i).conf.lowspeed     <= 'X';
        r.ch(i).conf.oddframe     <= 'X';
        r.ch(i).conf.interval     <= (others => '0');
        r.ch(i).conf.maxsize      <= (others => 'X');
        r.ch(i).conf.eptype       <= (others => 'X');
        r.ch(i).conf.address      <= (others => 'X');
        r.ch(i).conf.epnum        <= (others => 'X');

        r.ch(i).trans.epaddr      <= (others => '0');
        r.ch(i).trans.intervalcnt <= (others => '0');
        r.ch(i).trans.issued      <= '1';
        r.ch(i).trans.cnt         <= '0';
        r.ch(i).trans.seq         <= '0';
        r.ch(i).trans.size        <= (others => 'X');
        r.ch(i).trans.epaddr      <= (others => 'X');
        r.ch(i).trans.retries     <= (others => 'X');

        r.ch(i).intconf.datatogglerror           <= 'X';
        r.ch(i).intconf.crcerror                 <= 'X';
        r.ch(i).intconf.babble                   <= 'X';
        r.ch(i).intconf.transerror               <= 'X';
        r.ch(i).intconf.ack                      <= 'X';
        r.ch(i).intconf.nack                     <= 'X';
        r.ch(i).intconf.stall                    <= 'X';
        r.ch(i).intconf.cplt                     <= 'X';

        r.ch(i).intpend.datatogglerror           <= '0';
        r.ch(i).intpend.crcerror                 <= '0';
        r.ch(i).intpend.babble                   <= '0';
        r.ch(i).intpend.transerror               <= '0';
        r.ch(i).intpend.ack                      <= '0';
        r.ch(i).intpend.nack                     <= '0';
        r.ch(i).intpend.stall                    <= '0';
        r.ch(i).intpend.cplt                     <= '0';

      end loop;

    elsif rising_edge(usbclk_i) then
      r <= w;
    end if;
  end process;

  int_sync: entity work.sync
    generic map (
      RESET => '0'
    )
    port map (
      arst_i  => arst_i,
      clk_i   => clk_i,
      din_i   => int_s,
      dout_o  => int_sync_s
    );

  int_o <= int_sync_s;

  ahb2rdwr_inst: entity work.ahb2rdwr
    generic map (
      AWIDTH => 12, DWIDTH => 8
    )
    port map (
      clk_i     => usbclk_i,
      arst_i    => ausbrst_i,
      ahb_m2s_i => ahb_m2s_i,
      ahb_s2m_o => ahb_s2m_o,

      addr_o    => addr_s,
      dat_o     => dat_in_s,
      dat_i     => dat_out_s,
      rd_o      => rd_s,
      wr_o      => wr_s
    );


  hep_rd_s <= '1' when addr_s(10)='1' and rd_s='1' else '0' ;
  hep_wr_s <= '1' when addr_s(10)='1' and wr_s='1' else '0' ;

  epmem_inst: entity work.usb_epmem
    port map (
      uclk_i    => usbclk_i,
      urd_i     => epmem_read_en_s,
      uwr_i     => epmem_write_en_s,
      uaddr_i   => epmem_addr_s,
      udata_o   => epmem_data_out_s,
      udata_i   => epmem_data_in_s,

      hclk_i    => clk_i,
      hrd_i     => hep_rd_s,
      hwr_i     => hep_wr_s,
      haddr_i   => addr_s(9 downto 0),
      hdata_o   => hep_dat_s,
      hdata_i   => dat_in_s
  );

  usb_trans_inst: entity work.usb_trans
  port map (
    usbclk_i          => usbclk_i,
    ausbrst_i         => ausbrst_i,
    speed_i           => trans_speed_s,
    hostspeed_i       => r.speed,
    fs_ce_i           => fs_ce_s,
    usb_rst_i         => usb_rst_phy,
    -- Transmission
    pid_i             => trans_pid_s,

    -- Address/EP for token packets
    addr_i            => trans_addr_s,
    ep_i              => trans_ep_s,
    -- Frame number for SOF
    frame_i           => std_logic_vector(r.frame),
    --
    dsize_i           => trans_dsize_s,
    dsize_o           => trans_dsize_read_s,
    daddr_i           => trans_daddr_s,

    strobe_i          => trans_strobe_s,
    data_seq_i        => trans_data_seq_s,
    data_seq_valid_o  => trans_seq_valid_s,

    phy_txready_i     => Phy_TxReady,
    phy_txactive_i    => phy_txactive_s, -- from OE
    phy_txdata_o      => Phy_DataOut,
    phy_data_valid_o  => Phy_TxValid,
    phy_rxactive_i    => Phy_RxActive,
    phy_rxvalid_i     => Phy_RxValid,
    phy_rxdata_i      => Phy_DataIn,
    phy_rxerror_i     => Phy_RxError,
    phy_xcvrSelect_o  => Phy_XcvrSelect,

    -- Connection to EPMEM

    urd_o             => epmem_read_en_s,
    uwr_o             => epmem_write_en_s,
    uaddr_o           => epmem_addr_s,
    udata_i           => epmem_data_out_s,
    udata_o           => epmem_data_in_s,

    dbg_rx_data_done_o => dbg_rx_data_done_s,
    dbg_state_o        => dbg_trans_state_s,
    status_o            => trans_status_s,

    cnt_ack_o         =>  cnt_ack_s,
    cnt_nack_o        =>  cnt_nack_s,
    cnt_babble_o      =>  cnt_babble_s,
    cnt_stall_o       =>  cnt_stall_s ,
    cnt_crcerror_o    =>  cnt_crcerror_s,
    cnt_timeout_o     =>  cnt_timeout_s,
    cnt_errorpid_o    =>  cnt_errorpid_s,
    cnt_cplt_o        =>  cnt_cplt_s
  );

  process(usbclk_i)
  begin
    if rising_edge(usbclk_i) then
      read_data_r<=read_data_s;
    end if;
  end process;


  --epmem_addr_s <= std_logic_vector(r.epmem_addr);

  speed_o     <= r.speed;
  softcon_o   <= '0';
  noe_o       <= '0' when r.host_state=RESET1 else noe_s;
  vpo_o       <= '0' when r.host_state=RESET1 else vpo_s;
  vmo_o       <= '0' when r.host_state=RESET1 else vmo_s;
  int_async_o <= int_s;
  pwren_o     <= not r.sr.poweron;

  dat_out_s   <= hep_dat_s when addr_s(10)='1' else read_data_r;

  mode_o      <= '1';

  debubg: block
    signal fs: std_logic;
  begin
  debug: process(usbclk_i,ausbrst_i)
  begin
    if ausbrst_i='1' then
      dbg_o <= (others => '0');
      fs <= '0';
    elsif rising_edge(usbclk_i) then
        --dbg_o(0) <= Phy_RxActive;
        --dbg_o(1) <= Phy_TxActive_s;
        --dbg_o(2) <= fs;--Phy_RxError;
        --dbg_o(3) <= dbg_rx_data_done_s;--Phy_Linestate(0);
        --dbg_o(4) <= Phy_Linestate(1);

        --case r.host_state is
        --    when DETACHED | ATTACHED  => dbg_o(7 downto 5) <= "000";
        --    when IDLE                 => dbg_o(7 downto 5) <= "001";
        --    when RESET1 | RESET2      => dbg_o(7 downto 5) <= "010";
        --    when WAIT_SOF             => dbg_o(7 downto 5) <= "011";
        --    when IN1                  => dbg_o(7 downto 5) <= "100";
        --    when OUT1                 => dbg_o(7 downto 5) <= "101";
        --    when SOF1                 => dbg_o(7 downto 5) <= "110";
        --    when SETUP1               => dbg_o(7 downto 5) <= "111";
        --    when others               => dbg_o(7 downto 5) <= "111";
        --end case; 
        --
        --if fs_ce_s='1' then
        --  fs <= not fs;
        --end if;
        dbg_o(0) <= int_sync_s;
        dbg_o(1) <= r.intconfr.ginten;
        dbg_o(2) <= dbg_chan_interrupt_s(0);
        dbg_o(3) <= dbg_chan_interrupt_s(1);
        dbg_o(4) <= dbg_chan_interrupt_s(2);
    end if;
  end process;
  end block;
END rtl;

