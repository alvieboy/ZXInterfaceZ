entity SN74LCX245FT is
