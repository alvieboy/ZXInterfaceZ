library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity qspi is
  port (
    clk_i         : in std_logic;
    arst_i        : in std_logic;

  );
end entity qspi;

architecture beh of qspi is

begin

end architecture;

