
configuration t001 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t001);
        end for;
    end for;
end t001;

configuration t002 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t002);
        end for;
    end for;
end t002;

configuration t003 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t003);
        end for;
    end for;
end t003;

configuration t004 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t004);
        end for;
    end for;
end t004;

configuration t005 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t005);
        end for;
    end for;
end t005;

configuration t006 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t006);
        end for;
    end for;
end t006;

configuration t007 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t007);
        end for;
    end for;
end t007;

configuration t008 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t008);
        end for;
    end for;
end t008;

configuration t009 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t009);
        end for;
    end for;
end t009;

configuration t010 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t010);
        end for;
    end for;
end t010;

configuration t011 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t011);
        end for;
    end for;
end t011;

configuration t012 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t012);
        end for;
    end for;
end t012;

configuration t013 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t013);
        end for;
    end for;
end t013;

configuration t014 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t014);
        end for;
    end for;
end t014;

configuration t015 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t015);
        end for;
    end for;
end t015;

configuration t016 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t016);
        end for;
    end for;
end t016;

configuration t017 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t017);
        end for;
    end for;
end t017;

configuration t018 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t018);
        end for;
    end for;
end t018;


configuration t019 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t019);
        end for;
    end for;
end t019;

configuration t020 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t020);
        end for;
    end for;
end t020;

configuration t021 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t021);
        end for;
    end for;
end t021;
