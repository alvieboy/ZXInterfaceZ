
configuration t001 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t001);
        end for;
    end for;
end t001;

configuration t002 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t002);
        end for;
    end for;
end t002;

configuration t003 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t003);
        end for;
    end for;
end t003;

configuration t004 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t004);
        end for;
    end for;
end t004;

configuration t005 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t005);
        end for;
    end for;
end t005;

configuration t006 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t006);
        end for;
    end for;
end t006;

configuration t007 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t007);
        end for;
    end for;
end t007;
configuration t008 of tb_top is
    for sim
        for tbc: tbc_device
            use entity work.tbc_device(t008);
        end for;
    end for;
end t008;
